module m;
    // hello
    int a = 5 + 6;

    begin end
endmodule