initial 
	int a = 0;
