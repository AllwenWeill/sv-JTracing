module m;
    // hello
    int a = 5 + 6;
    int a;
    begin end
endmodule