module m;
    // hello
    int a = 5;

    begin end
endmodule