`include "file_defn.svh"
`define ID(x) x

module m;
    // hello
    string s = "FOO";

    begin end
endmodule

