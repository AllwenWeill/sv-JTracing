module m;
    // hello
    int a = 6 + 5;

    begin end
endmodule