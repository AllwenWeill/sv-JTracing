module m;
    // hello
    int a = 5 + 6;
    reg n;
    bit b;
    begin end
endmodule