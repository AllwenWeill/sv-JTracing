module m;
    // hello
    int a = 5 + 6;
    int n;
    begin end
endmodule