module m;
    // hello
    always_ff
    begin end
endmodule